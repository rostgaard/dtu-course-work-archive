--------------------------------------------------------------------------------
-- Wrapper other core generated DCM, to allow easy switching of the constants
--
-- Author     : Edgar Lakis <s081553@student.dtu.dk>
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.Vcomponents.all;

entity ClockDivider is
   generic(div : real);
   port(
      clkIn  : in  std_logic;
      clkOut : out std_logic
      );
end ClockDivider;



architecture DCM of ClockDivider is
begin
   -- use input clock, as no devision required
   copy_clock : if (div < 1.01) generate
      clkOut <= clkIn;
   end generate;

   -- divide the clock
   divide : if (div >= 1.01) generate
      alias CLKIN_IN  : std_logic is clkIn;
      alias CLKDV_OUT : std_logic is clkOut;

      signal CLKDV_BUF : std_logic;
      signal CLKFB_IN  : std_logic;
      signal CLK0_BUF  : std_logic;
      signal GND_BIT   : std_logic;
   begin
      --------------------------------------------------------------------------------
      -- Copyright (c) 1995-2008 Xilinx, Inc.  All rights reserved.
      --------------------------------------------------------------------------------
      --   ____  ____ 
      --  /   /\/   / 
      -- /___/  \  /    Vendor: Xilinx 
      -- \   \   \/     Version : 10.1.02
      --  \   \         Application : xaw2vhdl
      --  /   /         Filename : ClockDivider.vhd
      -- /___/   /\     Timestamp : 10/09/2009 12:40:50
      -- \   \  /  \ 
      --  \___\/\___\ 
      --
      --Command: xaw2vhdl-intstyle C:/Temp/actest/ClockDivider.xaw -st ClockDivider.vhd
      --Design Name:ClockDivider 
      --Device: xc2vp30-5ff896
      --
      -- Module ClockDivider 
      -- Generated by Xilinx Architecture Wizard
      -- Written for synthesis tool: XST

      GND_BIT <= '0';
      --   CLK0_OUT <= CLKFB_IN;
      CLKDV_BUFG_INST : BUFG
         port map (I => CLKDV_BUF,
                   O => CLKDV_OUT);

      CLK0_BUFG_INST : BUFG
         port map (I => CLK0_BUF,
                   O => CLKFB_IN);

      DCM_INST : DCM
         generic map(CLK_FEEDBACK          => "1X",
                     CLKDV_DIVIDE          => div,
                     CLKFX_DIVIDE          => 1,
                     CLKFX_MULTIPLY        => 4,
                     CLKIN_DIVIDE_BY_2     => false,
                     CLKIN_PERIOD          => 10.000,
                     CLKOUT_PHASE_SHIFT    => "NONE",
                     DESKEW_ADJUST         => "SYSTEM_SYNCHRONOUS",
                     DFS_FREQUENCY_MODE    => "LOW",
                     DLL_FREQUENCY_MODE    => "LOW",
                     DUTY_CYCLE_CORRECTION => true,
                     FACTORY_JF            => x"C080",
                     PHASE_SHIFT           => 0,
                     STARTUP_WAIT          => false)
         port map (CLKFB    => CLKFB_IN,
                   CLKIN    => CLKIN_IN,
                   DSSEN    => GND_BIT,
                   PSCLK    => GND_BIT,
                   PSEN     => GND_BIT,
                   PSINCDEC => GND_BIT,
                   RST      => GND_BIT,
                   CLKDV    => CLKDV_BUF,
                   CLKFX    => open,
                   CLKFX180 => open,
                   CLK0     => CLK0_BUF,
                   CLK2X    => open,
                   CLK2X180 => open,
                   CLK90    => open,
                   CLK180   => open,
                   CLK270   => open,
                   LOCKED   => open,
                   PSDONE   => open,
                   STATUS   => open);
   end generate;

end DCM;
