-- Listing 11.1
-- Single-port RAM with synchronous read
-- Modified from XST 8.1i rams_07
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity lc3_mem is
  generic(
    ADDR_WIDTH: integer:=12;
    DATA_WIDTH: integer:=8
    );
  port(
    clk: in std_logic;
	 reset: in std_logic;
	 rx: in std_logic;
	 tx: out std_logic;
    we, re: in std_logic; -- Write and read enable
    addr: in std_logic_vector(ADDR_WIDTH-1 downto 0);
    data: inout std_logic_vector(DATA_WIDTH-1 downto 0);
	 sw: in std_logic_vector(7 downto 0);
	 sseg_reg: out std_logic_vector(15 downto 0);
	 leds_reg: out std_logic_vector(7 downto 0);
	 btn: in std_logic_vector(4 downto 0)
    );
end lc3_mem;

architecture beh_arch of lc3_mem is
  type ram_type is array (0 to 2**ADDR_WIDTH-1)
    of std_logic_vector (DATA_WIDTH-1 downto 0);
  signal ram: ram_type := (
  -- Empty Traps/Interrupt Tables
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 0 - 7
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 8 - 15
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 16 - 23
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 24 - 31
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 32 - 39
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 40 - 47
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 48 - 55
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 56 - 63
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 64 - 71
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 72 - 79
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 80 - 87
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 88 - 95
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 96 - 103
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 104 - 111
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 112 - 119
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 120 - 127
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 128 - 135
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 136 - 143
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 144 - 151
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 152 - 159
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 160 - 167
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 168 - 175
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 176 - 183
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 184 - 191
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 192 - 199
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 200 - 207
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 208 - 215
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 216 - 223
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 224 - 231
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 232 - 239
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 240 - 247
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 248 - 255
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 256 - 263
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 264 - 271
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 272 - 279
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 280 - 287
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 288 - 295
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 296 - 303
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 304 - 311
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 312 - 319
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 320 - 327
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 328 - 335
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 336 - 343
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 344 - 351
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 352 - 359
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 360 - 367
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 368 - 375
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 376 - 383
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 384 - 391
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 392 - 399
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 400 - 407
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 408 - 415
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 416 - 423
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 424 - 431
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 432 - 439
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 440 - 447
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 448 - 455
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 456 - 463
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 464 - 471
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 472 - 479
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 480 - 487
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 488 - 495
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 496 - 503
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 504 - 511
-- Serial Port Program loader    (512-767)
X"2407", X"6080", X"07fe", X"6082", X"6284", X"07fe", X"7086", X"0ff9",  -- addr 512 - 519
X"fe00", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 520 - 527
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 528 - 535
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 536 - 543
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 544 - 551
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 552 - 559
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 560 - 567
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 568 - 575
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 576 - 583
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 584 - 591
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 592 - 599
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 600 - 607
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 608 - 615
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 616 - 623
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 624 - 631
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 632 - 639
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 640 - 647
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 648 - 655
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 656 - 663
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 664 - 671
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 672 - 679
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 680 - 687
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 688 - 695
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 696 - 703
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 704 - 711
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 712 - 719
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 720 - 727
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 728 - 735
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 736 - 743
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 744 - 751
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 752 - 759
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 760 - 767
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 768 - 775
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 776 - 783
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 784 - 791
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 792 - 799
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 800 - 807
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 808 - 815
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 816 - 823
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 824 - 831
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 832 - 839
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 840 - 847
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 848 - 855
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 856 - 863
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 864 - 871
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 872 - 879
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 880 - 887
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 888 - 895
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 896 - 903
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 904 - 911
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 912 - 919
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 920 - 927
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 928 - 935
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 936 - 943
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 944 - 951
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 952 - 959
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 960 - 967
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 968 - 975
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 976 - 983
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 984 - 991
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 992 - 999
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1000 - 1007
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1008 - 1015
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1016 - 1023
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1024 - 1031
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1032 - 1039
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1040 - 1047
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1048 - 1055
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1056 - 1063
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1064 - 1071
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1072 - 1079
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1080 - 1087
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1088 - 1095
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1096 - 1103
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1104 - 1111
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1112 - 1119
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1120 - 1127
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1128 - 1135
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1136 - 1143
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1144 - 1151
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1152 - 1159
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1160 - 1167
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1168 - 1175
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1176 - 1183
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1184 - 1191
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1192 - 1199
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1200 - 1207
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1208 - 1215
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1216 - 1223
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1224 - 1231
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1232 - 1239
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1240 - 1247
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1248 - 1255
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1256 - 1263
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1264 - 1271
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1272 - 1279
-- Start of user program         (1280-...)
X"2405", X"608a", X"7092", X"608e", X"7096", X"0ffb", X"fe00",  -- addr 1280 - 1286
 others => X"0000"
);
  signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);
  
  signal data_in: std_logic_vector(ADDR_WIDTH-1 downto 0);
  signal data_out: std_logic_vector(ADDR_WIDTH-1 downto 0);

  signal ram_signal: std_logic_vector(ADDR_WIDTH-1 downto 0);
  signal memory_map: std_logic_vector(ADDR_WIDTH-1 downto 0); 
  
  signal cs_mem: std_logic;
  
  signal cs_stdin_status: std_logic;
  signal cs_stdin_data: std_logic;
  
  signal cs_stdout_status: std_logic;
  signal cs_stdout_data: std_logic;
  
  signal cs_switch_data: std_logic;
  signal cs_btn_data: std_logic;
  signal cs_sseg: std_logic;
  signal cs_led: std_logic;
  
  --uart specific
  signal uart_w_data: std_logic_vector(7 downto 0);
  signal uart_r_data: std_logic_vector(7 downto 0);
  signal tx_full, rx_empty: std_logic;
  
begin

   -- instantiate uart
   uart_unit: entity work.uart(str_arch)
      port map(clk=>clk, 
					reset=>reset, 
					rd_uart=> cs_stdin_status,
               wr_uart=> cs_stdout_status,
					rx=>rx, 
					w_data=>uart_w_data,
               tx_full=>tx_full, 
					rx_empty=>rx_empty,
               r_data=>uart_r_data, 
					tx=>tx);



  process (addr_reg)
  begin
    cs_mem <= '0';
	 cs_stdin_status <= '0';
	 cs_stdin_data <= '0';
	 cs_stdout_status <= '0';
	 cs_stdout_data <= '0';
	 cs_switch_data <= '0';
	 cs_btn_data <= '0';
	 cs_sseg <= '0';
	 cs_led <= '0';
   
	 if addr_reg >= X"0000" AND addr_reg <= X"DFFF" then --reserved space in software memory, rest is for I/O
	   cs_mem <= '1';
		-- xFE00 Stdin Status Register
    elsif addr_reg = X"FE00" then
	   cs_stdin_status <= '1';
		-- xFE02 Stdin Data Register
    elsif addr_reg = X"FE02" then
		cs_stdin_data <= '1';
		-- xFE04 Stdout Status Register
	 elsif addr_reg = X"FE04" then
		cs_stdout_status <= '1';
		 -- xFE06 Stdout Data Register
	 elsif addr_reg = X"FE06" then
		cs_stdout_data <= '1';
		-- xFE0A Switches Data Register
	 elsif addr_reg = X"FE0A" then
		cs_switch_data <= '1';
		-- xFE0E Buttons Data Register
	 elsif addr_reg = X"FE0E" then
		cs_btn_data <= '1';
		-- xFE12 7SegDisplay Data Register
	 elsif addr_reg = X"FE12" then
		cs_sseg <= '1';
		 -- xFE16 Leds Data Register
	 elsif addr_reg = X"FE16" then
		cs_led <= '1';
    end if;
  end process;
 
  -- RAM template
  --data <= ram(to_integer(unsigned(addr_reg))) when re = '1' and cs_mem = '1' 
    --else (others => 'Z');
  
  --process (clk)
  --begin
    --if (clk'event and clk = '1') then
     --if (we='1') and cs_mem = '1' then
       --ram(to_integer(unsigned(addr))) <= data;
     --end if;
    -- addr_reg <= addr;
   --end if;
 -- end process;
  
  	-- cs_mem is In/Out
  data <= ram(to_integer(unsigned(addr_reg))) when re = '1' and cs_mem = '1' 
    else (others => 'Z');
	 
  process (clk)
  begin
    if (clk'event and clk = '1') then
      if (we='1') and cs_stdin_status = '1' then
        ram(to_integer(unsigned(addr))) <= data;
      end if;
      addr_reg <= addr;
    end if;
  end process;
  
	-- cs_stdin_status is out
  data <= not rx_empty & "000" & X"000" when re = '1' and cs_stdin_status = '1' 
    else (others => 'Z');
  
	-- cs_stdin_data  is out
  data <= uart_r_data when re = '1' and cs_stdin_data = '1' 
    else (others => 'Z');
  
	-- cs_stdout_status  is out
  data <= not tx_full & "000" & X"000" when re = '1' and cs_stdout_status = '1' 
    else (others => 'Z');
	 
	-- cs_stout_data is in 
  process (clk)
  begin
    if (clk'event and clk = '1') then
      if (we='1') and cs_stdout_data = '1' then
        uart_w_data <= data;
      end if;
    end if;
  end process;
  
  --cs_switch_data  is out
  data <= sw when re = '1' and cs_switch_data = '1' 
    else (others => 'Z');
	 
  -- TODO cs_btn_data  is out
  data <= X"00" & "000" & btn when re = '1' and cs_btn_data = '1' 
    else (others => 'Z');
	 
	-- cs_sseg  is in 
  process (clk)
  begin
    if (clk'event and clk = '1') then
      if (we='1') and cs_sseg = '1' then
        sseg_reg <= data;
      end if;
    end if;
  end process;
  
 	-- cs_leds  is in 
  process (clk)
  begin
    if (clk'event and clk = '1') then
      if (we='1') and cs_led = '1' then
        leds_reg <= data;
      end if;
    end if;
  end process;
        
end beh_arch;
