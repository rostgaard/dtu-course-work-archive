----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:20:39 02/26/2010 
-- Design Name: 
-- Module Name:    reg_reset - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.ALL;
 
entity reg_reset is
	port(
		clk,reset: in std_logic;
		d: in std_logic_vector(7 downto 0);
		q: out std_logic_vector(7 downto 0)
	);
end reg_reset;

architecture arch of reg_reset is
begin 
	process(clk,reset)
	begin
		if (reset='1') then
			q <=(others => '0');
		elsif (clk'event and clk = '1') then
			q <= d;
		end if;
	end process;
end arch;