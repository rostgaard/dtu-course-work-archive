-- Listing 11.1
-- Single-port RAM with synchronous read
-- Modified from XST 8.1i rams_07
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity lc3_mem is
  generic(
    ADDR_WIDTH: integer:=12;
    DATA_WIDTH: integer:=8
    );
  port(
    clk: in std_logic;
	 reset: in std_logic;
	 rx: in std_logic;
	 tx: out std_logic;
    we, re: in std_logic; -- Write and read enable
    addr: in std_logic_vector(ADDR_WIDTH-1 downto 0);
    data: inout std_logic_vector(DATA_WIDTH-1 downto 0);
	 sw: in std_logic_vector(7 downto 0);
	 sseg_reg: out std_logic_vector(15 downto 0);
	 leds_reg: out std_logic_vector(7 downto 0);
	 btn: in std_logic_vector(4 downto 0)
    );
end lc3_mem;

architecture beh_arch of lc3_mem is
  type ram_type is array (0 to 2**ADDR_WIDTH-1)
    of std_logic_vector (DATA_WIDTH-1 downto 0);
  signal ram: ram_type := (
-- Trap Vector Table             (0-255)
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 0 - 7
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 8 - 15
X"0349", X"0349", X"0358", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 16 - 23
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 24 - 31
X"035a", X"035e", X"0364", X"0371", X"037d", X"0300", X"0349", X"0349",  -- addr 32 - 39
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 40 - 47
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 48 - 55
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 56 - 63
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 64 - 71
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 72 - 79
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 80 - 87
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 88 - 95
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 96 - 103
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 104 - 111
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 112 - 119
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 120 - 127
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 128 - 135
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 136 - 143
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 144 - 151
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 152 - 159
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 160 - 167
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 168 - 175
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 176 - 183
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 184 - 191
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 192 - 199
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 200 - 207
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 208 - 215
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 216 - 223
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 224 - 231
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 232 - 239
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 240 - 247
X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349", X"0349",  -- addr 248 - 255
-- Interrupt Vector Table        (256-511)
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 256 - 263
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 264 - 271
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 272 - 279
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 280 - 287
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 288 - 295
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 296 - 303
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 304 - 311
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 312 - 319
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 320 - 327
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 328 - 335
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 336 - 343
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 344 - 351
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 352 - 359
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 360 - 367
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 368 - 375
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 376 - 383
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 384 - 391
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 392 - 399
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 400 - 407
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 408 - 415
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 416 - 423
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 424 - 431
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 432 - 439
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 440 - 447
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 448 - 455
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 456 - 463
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 464 - 471
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 472 - 479
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 480 - 487
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 488 - 495
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"034f",  -- addr 496 - 503
X"034f", X"034f", X"034f", X"034f", X"034f", X"034f", X"0352", X"0355",  -- addr 504 - 511
-- Serial Port Program loader    (512-767)
X"e00b", X"48c4", X"2007", X"b003", X"2006", X"b002", X"0e26", X"fe16",  -- addr 512 - 519
X"fe12", X"fe00", X"00ff", X"cccc", X"000a", X"002d", X"002d", X"002d",  -- addr 520 - 527
X"0020", X"0057", X"0061", X"0069", X"0074", X"0069", X"006e", X"0067",  -- addr 528 - 535
X"0020", X"0066", X"006f", X"0072", X"0020", X"0070", X"0072", X"006f",  -- addr 536 - 543
X"0067", X"0072", X"0061", X"006d", X"002e", X"002e", X"002e", X"000a",  -- addr 544 - 551
X"0000", X"ffe5", X"ffaf", X"ffab", X"ffad", X"48a1", X"23fa", X"1001",  -- addr 552 - 559
X"0bfc", X"489d", X"23f7", X"1201", X"0407", X"23f5", X"1201", X"040e",  -- addr 560 - 567
X"23f3", X"1201", X"046a", X"0ff1", X"e002", X"4888", X"0fee", X"0052",  -- addr 568 - 575
X"0065", X"0061", X"0064", X"0079", X"002e", X"0000", X"488e", X"1820",  -- addr 576 - 583
X"b1bf", X"488b", X"1a20", X"b1bc", X"4888", X"bbba", X"7140", X"1b61",  -- addr 584 - 591
X"193f", X"03fa", X"e002", X"4872", X"0fd8", X"000a", X"0050", X"0072",  -- addr 592 - 599
X"006f", X"0067", X"0072", X"0061", X"006d", X"006d", X"0069", X"006e",  -- addr 600 - 607
X"0067", X"0020", X"0064", X"006f", X"006e", X"0065", X"002e", X"000a",  -- addr 608 - 615
X"002d", X"002d", X"002d", X"0020", X"0050", X"0072", X"0065", X"0073",  -- addr 616 - 623
X"0073", X"0020", X"0072", X"0065", X"0073", X"0065", X"0074", X"0028",  -- addr 624 - 631
X"0045", X"004e", X"0054", X"0045", X"0052", X"0020", X"0070", X"0075",  -- addr 632 - 639
X"0073", X"0068", X"002d", X"0062", X"0075", X"0074", X"0074", X"006f",  -- addr 640 - 647
X"006e", X"0029", X"0020", X"006f", X"0072", X"0020", X"0070", X"0072",  -- addr 648 - 655
X"006f", X"0067", X"0072", X"0061", X"006d", X"0020", X"006e", X"0065",  -- addr 656 - 663
X"0078", X"0074", X"0020", X"0062", X"006c", X"006f", X"0063", X"006b",  -- addr 664 - 671
X"002e", X"002e", X"002e", X"000a", X"0000", X"5020", X"b160", X"b160",  -- addr 672 - 679
X"e003", X"481c", X"482a", X"c000", X"000a", X"004a", X"0075", X"006d",  -- addr 680 - 687
X"0070", X"0069", X"006e", X"0067", X"0020", X"0074", X"006f", X"0020",  -- addr 688 - 695
X"0075", X"0073", X"0065", X"0072", X"0020", X"0063", X"006f", X"0064",  -- addr 696 - 703
X"0065", X"002e", X"000a", X"0000", X"fe04", X"fe06", X"1220", X"6040",  -- addr 704 - 711
X"0405", X"a5fa", X"07fe", X"b1f9", X"1261", X"0ff9", X"c1c0", X"2539",  -- addr 712 - 719
X"6080", X"07fe", X"6082", X"c1c0", X"0100", X"2533", X"6080", X"07fe",  -- addr 720 - 727
X"6082", X"6280", X"07fe", X"6282", X"25f7", X"1080", X"1000", X"07fe",  -- addr 728 - 735
X"1000", X"1040", X"c1c0", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 736 - 743
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 744 - 751
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 752 - 759
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 760 - 767
-- Trap Implementation           (768-1279)
X"e006", X"f022", X"a09d", X"229f", X"5001", X"b09a", X"c1c0", X"000a",  -- addr 768 - 775
X"000a", X"002d", X"002d", X"002d", X"0020", X"0068", X"0061", X"006c",  -- addr 776 - 783
X"0074", X"0069", X"006e", X"0067", X"0020", X"0074", X"0068", X"0065",  -- addr 784 - 791
X"0020", X"004c", X"0043", X"002d", X"0033", X"0020", X"002d", X"002d",  -- addr 792 - 799
X"002d", X"000a", X"000a", X"0000", X"000a", X"000a", X"002d", X"002d",  -- addr 800 - 807
X"002d", X"0020", X"0075", X"006e", X"0064", X"0065", X"0066", X"0069",  -- addr 808 - 815
X"006e", X"0065", X"0064", X"0020", X"0074", X"0072", X"0061", X"0070",  -- addr 816 - 823
X"0020", X"0065", X"0078", X"0065", X"0063", X"0075", X"0074", X"0065",  -- addr 824 - 831
X"0064", X"0020", X"002d", X"002d", X"002d", X"000a", X"000a", X"0000",  -- addr 832 - 839
X"eeee", X"21fe", X"b057", X"0fb4", X"e1d7", X"f022", X"0fb1", X"5020",  -- addr 840 - 847
X"103d", X"0ff8", X"5020", X"103e", X"0ff5", X"5020", X"103f", X"0ff2",  -- addr 848 - 855
X"b049", X"c1c0", X"a041", X"07fe", X"a040", X"c1c0", X"3246", X"a23e",  -- addr 856 - 863
X"07fe", X"b03d", X"2242", X"c1c0", X"3042", X"3242", X"3e44", X"1220",  -- addr 864 - 871
X"6040", X"0403", X"f021", X"1261", X"0ffb", X"2039", X"2239", X"2e3b",  -- addr 872 - 879
X"c1c0", X"3e34", X"e039", X"f022", X"f020", X"f021", X"3030", X"5020",  -- addr 880 - 887
X"102a", X"f021", X"202c", X"2e2a", X"c1c0", X"3029", X"3229", X"3429",  -- addr 888 - 895
X"3629", X"3e29", X"1220", X"6440", X"201f", X"5002", X"040f", X"f021",  -- addr 896 - 903
X"5020", X"1628", X"1000", X"14a0", X"0601", X"1021", X"1482", X"16ff",  -- addr 904 - 911
X"03f9", X"1020", X"0403", X"f021", X"1261", X"0fed", X"2010", X"2210",  -- addr 912 - 919
X"2410", X"2610", X"2e10", X"c1c0", X"fe00", X"fe02", X"fe04", X"fe06",  -- addr 920 - 927
X"fffe", X"fe10", X"fe12", X"7fff", X"00ff", X"0000", X"0000", X"0000",  -- addr 928 - 935
X"0000", X"0000", X"0000", X"0000", X"000a", X"0049", X"006e", X"0070",  -- addr 936 - 943
X"0075", X"0074", X"0020", X"0061", X"0020", X"0063", X"0068", X"0061",  -- addr 944 - 951
X"0072", X"0061", X"0063", X"0074", X"0065", X"0072", X"003e", X"0020",  -- addr 952 - 959
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 960 - 967
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 968 - 975
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 976 - 983
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 984 - 991
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 992 - 999
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1000 - 1007
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1008 - 1015
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1016 - 1023
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1024 - 1031
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1032 - 1039
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1040 - 1047
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1048 - 1055
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1056 - 1063
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1064 - 1071
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1072 - 1079
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1080 - 1087
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1088 - 1095
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1096 - 1103
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1104 - 1111
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1112 - 1119
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1120 - 1127
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1128 - 1135
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1136 - 1143
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1144 - 1151
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1152 - 1159
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1160 - 1167
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1168 - 1175
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1176 - 1183
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1184 - 1191
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1192 - 1199
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1200 - 1207
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1208 - 1215
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1216 - 1223
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1224 - 1231
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1232 - 1239
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1240 - 1247
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1248 - 1255
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1256 - 1263
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1264 - 1271
X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  -- addr 1272 - 1279
-- Start of user program         (1280-...)
X"e004", X"f022", X"2001", X"c000", X"0916", X"000a", X"0020", X"002a",  -- addr 1280 - 1287
X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a",  -- addr 1288 - 1295
X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a",  -- addr 1296 - 1303
X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a",  -- addr 1304 - 1311
X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a",  -- addr 1312 - 1319
X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a",  -- addr 1320 - 1327
X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a",  -- addr 1328 - 1335
X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a",  -- addr 1336 - 1343
X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a",  -- addr 1344 - 1351
X"002a", X"000a", X"0020", X"002a", X"0020", X"0020", X"0054", X"0068",  -- addr 1352 - 1359
X"0069", X"0073", X"0020", X"0075", X"0073", X"0065", X"0072", X"0020",  -- addr 1360 - 1367
X"0070", X"0072", X"006f", X"0067", X"0072", X"0061", X"006d", X"0020",  -- addr 1368 - 1375
X"0064", X"006f", X"0065", X"0073", X"006e", X"0027", X"0074", X"0020",  -- addr 1376 - 1383
X"0064", X"006f", X"0020", X"0061", X"006e", X"0079", X"0074", X"0068",  -- addr 1384 - 1391
X"0069", X"006e", X"0067", X"0020", X"0069", X"006e", X"0074", X"0065",  -- addr 1392 - 1399
X"0072", X"0065", X"0073", X"0074", X"0069", X"006e", X"0067", X"002e",  -- addr 1400 - 1407
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1408 - 1415
X"0020", X"0020", X"0020", X"0020", X"002a", X"000a", X"0020", X"002a",  -- addr 1416 - 1423
X"0020", X"0020", X"0059", X"006f", X"0075", X"0020", X"0073", X"0068",  -- addr 1424 - 1431
X"006f", X"0075", X"006c", X"0064", X"0020", X"0074", X"0072", X"0079",  -- addr 1432 - 1439
X"0020", X"0074", X"006f", X"0020", X"0075", X"0070", X"006c", X"006f",  -- addr 1440 - 1447
X"0061", X"0064", X"0020", X"0079", X"006f", X"0075", X"0072", X"0020",  -- addr 1448 - 1455
X"006f", X"0077", X"006e", X"0020", X"0070", X"0072", X"006f", X"0067",  -- addr 1456 - 1463
X"0072", X"0061", X"006d", X"003a", X"0020", X"0020", X"0020", X"0020",  -- addr 1464 - 1471
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1472 - 1479
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1480 - 1487
X"002a", X"000a", X"0020", X"002a", X"0020", X"0020", X"0020", X"0020",  -- addr 1488 - 1495
X"0031", X"002e", X"0020", X"0043", X"006f", X"006d", X"0070", X"0069",  -- addr 1496 - 1503
X"006c", X"0065", X"0020", X"0079", X"006f", X"0075", X"0072", X"0020",  -- addr 1504 - 1511
X"0070", X"0072", X"006f", X"0067", X"0072", X"0061", X"006d", X"0020",  -- addr 1512 - 1519
X"0028", X"0070", X"0072", X"006f", X"0064", X"0075", X"0063", X"0065",  -- addr 1520 - 1527
X"0020", X"002e", X"006f", X"0062", X"006a", X"0020", X"0066", X"0069",  -- addr 1528 - 1535
X"006c", X"0065", X"0029", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1536 - 1543
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1544 - 1551
X"0020", X"0020", X"0020", X"0020", X"002a", X"000a", X"0020", X"002a",  -- addr 1552 - 1559
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"005b",  -- addr 1560 - 1567
X"006f", X"0070", X"0074", X"0069", X"006f", X"006e", X"0031", X"005d",  -- addr 1568 - 1575
X"0020", X"0055", X"0073", X"0065", X"0020", X"004c", X"0043", X"0033",  -- addr 1576 - 1583
X"0045", X"0064", X"0069", X"0074", X"002e", X"0065", X"0078", X"0065",  -- addr 1584 - 1591
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1592 - 1599
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1600 - 1607
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1608 - 1615
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1616 - 1623
X"002a", X"000a", X"0020", X"002a", X"0020", X"0020", X"0020", X"0020",  -- addr 1624 - 1631
X"0020", X"0020", X"0020", X"005b", X"006f", X"0070", X"0074", X"0069",  -- addr 1632 - 1639
X"006f", X"006e", X"0032", X"005d", X"0020", X"0055", X"0073", X"0065",  -- addr 1640 - 1647
X"0020", X"004c", X"0043", X"0033", X"0020", X"0063", X"006f", X"006d",  -- addr 1648 - 1655
X"006d", X"0061", X"006e", X"0064", X"0020", X"006c", X"0069", X"006e",  -- addr 1656 - 1663
X"0065", X"0020", X"0061", X"0073", X"0073", X"0065", X"006d", X"0062",  -- addr 1664 - 1671
X"006c", X"0065", X"0072", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1672 - 1679
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1680 - 1687
X"0020", X"0020", X"0020", X"0020", X"002a", X"000a", X"0020", X"002a",  -- addr 1688 - 1695
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1696 - 1703
X"0020", X"0020", X"006c", X"0063", X"0033", X"0061", X"0073", X"0020",  -- addr 1704 - 1711
X"0061", X"0073", X"006d", X"005f", X"0073", X"006f", X"0075", X"0072",  -- addr 1712 - 1719
X"0063", X"0065", X"002e", X"0061", X"0073", X"006d", X"0020", X"0020",  -- addr 1720 - 1727
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1728 - 1735
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1736 - 1743
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1744 - 1751
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1752 - 1759
X"002a", X"000a", X"0020", X"002a", X"0020", X"0020", X"0020", X"0020",  -- addr 1760 - 1767
X"0020", X"0020", X"0020", X"005b", X"006f", X"0070", X"0074", X"0069",  -- addr 1768 - 1775
X"006f", X"006e", X"0033", X"005d", X"0020", X"0043", X"006f", X"006d",  -- addr 1776 - 1783
X"0070", X"0069", X"006c", X"0065", X"0020", X"0043", X"0020", X"0073",  -- addr 1784 - 1791
X"006f", X"0075", X"0072", X"0063", X"0065", X"0020", X"0020", X"0020",  -- addr 1792 - 1799
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1800 - 1807
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1808 - 1815
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1816 - 1823
X"0020", X"0020", X"0020", X"0020", X"002a", X"000a", X"0020", X"002a",  -- addr 1824 - 1831
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1832 - 1839
X"0020", X"0020", X"006c", X"0063", X"0063", X"0020", X"002d", X"006f",  -- addr 1840 - 1847
X"0020", X"0063", X"005f", X"0073", X"006f", X"0075", X"0072", X"0063",  -- addr 1848 - 1855
X"0065", X"002e", X"006f", X"0062", X"006a", X"0020", X"0063", X"005f",  -- addr 1856 - 1863
X"0073", X"006f", X"0075", X"0072", X"0063", X"0065", X"002e", X"0063",  -- addr 1864 - 1871
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1872 - 1879
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1880 - 1887
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 1888 - 1895
X"002a", X"000a", X"0020", X"002a", X"0020", X"0020", X"0020", X"0020",  -- addr 1896 - 1903
X"0032", X"002e", X"0020", X"0041", X"0063", X"0074", X"0069", X"0076",  -- addr 1904 - 1911
X"0061", X"0074", X"0065", X"0020", X"0070", X"0072", X"006f", X"0067",  -- addr 1912 - 1919
X"0072", X"0061", X"006d", X"006d", X"0065", X"0072", X"0020", X"006f",  -- addr 1920 - 1927
X"006e", X"0020", X"0046", X"0050", X"0047", X"0041", X"0020", X"0028",  -- addr 1928 - 1935
X"0070", X"0075", X"0073", X"0068", X"0020", X"0060", X"004c", X"0045",  -- addr 1936 - 1943
X"0046", X"0054", X"0027", X"0020", X"0070", X"0075", X"0073", X"0068",  -- addr 1944 - 1951
X"002d", X"0062", X"0075", X"0074", X"0074", X"006f", X"006e", X"0029",  -- addr 1952 - 1959
X"0020", X"0020", X"0020", X"0020", X"002a", X"000a", X"0020", X"002a",  -- addr 1960 - 1967
X"0020", X"0020", X"0020", X"0020", X"0033", X"002e", X"0020", X"0052",  -- addr 1968 - 1975
X"0069", X"0067", X"0068", X"0074", X"0020", X"0063", X"006c", X"0069",  -- addr 1976 - 1983
X"0063", X"006b", X"0020", X"006f", X"006e", X"0020", X"002e", X"006f",  -- addr 1984 - 1991
X"0062", X"006a", X"0020", X"0066", X"0069", X"006c", X"0065", X"0020",  -- addr 1992 - 1999
X"0061", X"006e", X"0064", X"0020", X"0073", X"0065", X"006c", X"0065",  -- addr 2000 - 2007
X"0063", X"0074", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 2008 - 2015
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 2016 - 2023
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 2024 - 2031
X"002a", X"000a", X"0020", X"002a", X"0020", X"0020", X"0020", X"0020",  -- addr 2032 - 2039
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0043", X"003a",  -- addr 2040 - 2047
X"005c", X"006c", X"0063", X"0033", X"005c", X"0062", X"0069", X"006e",  -- addr 2048 - 2055
X"005c", X"004c", X"0043", X"0033", X"0054", X"0065", X"0072", X"006d",  -- addr 2056 - 2063
X"0069", X"006e", X"0061", X"006c", X"002e", X"0065", X"0078", X"0065",  -- addr 2064 - 2071
X"0020", X"0069", X"006e", X"0020", X"0022", X"004f", X"0070", X"0065",  -- addr 2072 - 2079
X"006e", X"0020", X"0077", X"0069", X"0074", X"0068", X"0022", X"0020",  -- addr 2080 - 2087
X"0064", X"0069", X"0061", X"006c", X"006f", X"0067", X"0020", X"0020",  -- addr 2088 - 2095
X"0020", X"0020", X"0020", X"0020", X"002a", X"000a", X"0020", X"002a",  -- addr 2096 - 2103
X"0020", X"0020", X"0020", X"0020", X"0034", X"002e", X"0020", X"0057",  -- addr 2104 - 2111
X"0061", X"0069", X"0074", X"0020", X"0066", X"006f", X"0072", X"0020",  -- addr 2112 - 2119
X"0070", X"0072", X"006f", X"0067", X"0072", X"0061", X"006d", X"006d",  -- addr 2120 - 2127
X"0069", X"006e", X"0067", X"0020", X"0074", X"006f", X"0020", X"0066",  -- addr 2128 - 2135
X"0069", X"006e", X"0069", X"0073", X"0068", X"0020", X"0020", X"0020",  -- addr 2136 - 2143
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 2144 - 2151
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 2152 - 2159
X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020", X"0020",  -- addr 2160 - 2167
X"002a", X"000a", X"0020", X"002a", X"0020", X"0020", X"0020", X"0020",  -- addr 2168 - 2175
X"0020", X"0020", X"0020", X"0054", X"0068", X"0065", X"0020", X"0049",  -- addr 2176 - 2183
X"002f", X"004f", X"0020", X"0062", X"006f", X"0061", X"0072", X"0064",  -- addr 2184 - 2191
X"0020", X"006c", X"0065", X"0064", X"0073", X"0020", X"0077", X"0069",  -- addr 2192 - 2199
X"006c", X"006c", X"0020", X"0067", X"006f", X"0020", X"006f", X"0066",  -- addr 2200 - 2207
X"0066", X"0020", X"0061", X"006e", X"0064", X"0020", X"006d", X"0065",  -- addr 2208 - 2215
X"0073", X"0073", X"0061", X"0067", X"0065", X"0020", X"0077", X"0069",  -- addr 2216 - 2223
X"006c", X"006c", X"0020", X"0061", X"0070", X"0070", X"0065", X"0061",  -- addr 2224 - 2231
X"0072", X"002e", X"0020", X"0020", X"002a", X"000a", X"0020", X"002a",  -- addr 2232 - 2239
X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a",  -- addr 2240 - 2247
X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a",  -- addr 2248 - 2255
X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a",  -- addr 2256 - 2263
X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a",  -- addr 2264 - 2271
X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a",  -- addr 2272 - 2279
X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a",  -- addr 2280 - 2287
X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a",  -- addr 2288 - 2295
X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a", X"002a",  -- addr 2296 - 2303
X"002a", X"000a", X"000a", X"0000", X"004b", X"0065", X"0079", X"0020",  -- addr 2304 - 2311
X"0070", X"0072", X"0065", X"0073", X"0073", X"0065", X"0064", X"003a",  -- addr 2312 - 2319
X"0020", X"005b", X"0020", X"005d", X"000a", X"0000", X"e3ed", X"e5fe",  -- addr 2320 - 2327
X"14bc", X"f020", X"7080", X"1060", X"f022", X"0ffb",  -- addr 2328 - 2333
others => X"0000"

);
  signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);

  -- Chip selector signals
  signal cs_mem: std_logic;
  signal cs_stdin_status: std_logic;
  signal uart_rd_en: std_logic;
  signal cs_stdout_status: std_logic;
  signal uart_wr_en: std_logic;
  signal cs_switch_data: std_logic;
  signal cs_btn_data: std_logic;
  signal cs_sseg: std_logic;
  signal cs_led: std_logic;
  
  -- uart specific signals
  signal uart_w_data: std_logic_vector(7 downto 0);
  signal uart_r_data: std_logic_vector(7 downto 0);
  signal tx_full, rx_empty: std_logic;
  
begin

   -- instantiate uart
   uart_unit: entity work.uart(str_arch)
      port map(clk=>clk, 
					reset=>reset, 
					rd_uart=> uart_rd_en,
               wr_uart=> uart_wr_en,
					rx=>rx, 
					w_data=>uart_w_data,
               tx_full=>tx_full, 
					rx_empty=>rx_empty,
               r_data=>uart_r_data, 
					tx=>tx);

  --reserved space in software memory, rest is for I/O
	cs_mem <= '1' when addr >= X"0000" and addr <= X"DFFF" else '0';
  -- cs_mem is In/Out. This is the main memory
  data <= ram(to_integer(unsigned(addr_reg))) when re = '1' and cs_mem = '1' 
    else (others => 'Z');
	 
  process (clk)
  begin
    if (clk'event and clk = '1') then
      if (we='1') and cs_mem = '1' then
        ram(to_integer(unsigned(addr))) <= data;
      end if;
      addr_reg <= addr;
    end if;
  end process;


  -- xFE00 Stdin Status Register
  cs_stdin_status <= '1' when addr = X"FE00" and re = '1' else '0';
  data <= not rx_empty & "000" & X"000" when cs_stdin_status = '1' 
    else (others => 'Z');

  -- xFE02 Stdin Data Register, uart_rd_en acts as chip select
  uart_rd_en <= '1' when addr = X"FE02" and re = '1' else '0';
	-- cs_stdin_data  is out
  data <= uart_r_data when uart_rd_en = '1' 
    else (others => 'Z');

  -- xFE04 Stdout Status Register
  cs_stdout_status <= '1' when re = '1' and addr = X"FE04" else '0';
	-- cs_stdout_status  is out
  data <= not tx_full & "000" & X"000" when cs_stdout_status = '1' 
    else (others => 'Z');		

  -- xFE06 Stdout Data Register
  uart_wr_en <= '1' when addr = X"FE06" and we = '1' else '0';
 	-- cs_stout_data is in 
  uart_w_data <= data(7 downto 0);

  -- xFE0A Switches Data Register
  cs_switch_data <= '1' when addr = X"FE0A" and re = '1' else '0';
  --cs_switch_data  is out
  data <= sw when re = '1' and cs_switch_data = '1' 
    else (others => 'Z');		

  -- xFE0E Buttons Data Register
  cs_btn_data <= '1' when addr = X"FE0E" and re = '1' else '0';
  -- cs_btn_data  is out
  data <= X"00" & "000" & btn when cs_btn_data = '1' 
    else (others => 'Z');

  -- xFE12 7SegDisplay Data Register
  cs_sseg <= '1' when addr = X"FE12" and we='1' else '0';
	-- cs_sseg  is in 
  process (clk)
  begin
    if (clk'event and clk = '1') then
      if cs_sseg = '1' then
        sseg_reg <= data;
      end if;
    end if;
  end process;		

  -- xFE16 Leds Data Register
  cs_led <= '1' when addr = X"FE16" and we='1' else '0';
 	-- cs_leds  is in 
  process (clk)
  begin
    if (clk'event and clk = '1') then
      if cs_led = '1' then
        leds_reg <= data (7 downto 0);
      end if;
    end if;
  end process;
      
end beh_arch;
